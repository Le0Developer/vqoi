module vqoi

pub struct Image {
pub:
	pixels [][4]byte
	metadata ImageMetadata
}
