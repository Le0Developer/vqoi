module vqoi

pub struct Image {
pub:
	rgba [][4]byte
	metadata ImageMetadata
}
