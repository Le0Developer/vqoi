module vqoi

pub struct Image {
pub:
	rgba [][4]u8
	metadata ImageMetadata
}
